module LR_Keymill(clk, rst, key, load_key, iv, load_iv, run, stream_out, output_ready);
	input clk, rst, load_key, load_iv, run;
	input [7:0] key, iv;
	output output_ready;
	output [7:0] stream_out;
	reg output_ready;
	reg [7:0] stream_out;
	
	reg [0:30] R1;
	reg [0:31] R2, R3;
	reg [0:32] R4;
	
	reg [2:0] ready_counter;
	reg warm_up_done;
	
	wire F1p1_, F2p1_, F3p1_, F4p1_, F1p1, F2p1, F3p1, F4p1;
	wire F1p2_, F2p2_, F3p2_, F4p2_, F1p2, F2p2, F3p2, F4p2;
	wire F1p3_, F2p3_, F3p3_, F4p3_, F1p3, F2p3, F3p3, F4p3;
	wire F1p4_, F2p4_, F3p4_, F4p4_, F1p4, F2p4, F3p4, F4p4;
	wire F1p5_, F2p5_, F3p5_, F4p5_, F1p5, F2p5, F3p5, F4p5;
	wire F1p6_, F2p6_, F3p6_, F4p6_, F1p6, F2p6, F3p6, F4p6;
	wire F1p7_, F2p7_, F3p7_, F4p7_, F1p7, F2p7, F3p7, F4p7;
	wire F1p8_, F2p8_, F3p8_, F4p8_, F1p8, F2p8, F3p8, F4p8;
	
	reg [2:0] state;
	parameter State_RST = 3'b000, State_Load_Key = 3'b001, State_Load_IV = 3'b010, State_Warm_Up = 3'b011, State_Gen_Output=3'b100, State_Halt=3'b101;
	
	always @(posedge clk or negedge rst)
		if (~rst)
			state <= State_RST;
		else
			case (state)
			State_RST: begin
				stream_out <= 1'b0;
				output_ready <= 1'b0;
				ready_counter <= 3'b000;
				warm_up_done <= 1'b0;
				
				if (load_key)
					state <= State_Load_Key;
				else
					state <= State_RST;
				end
			
			State_Load_Key: begin		
					R1[23:30] <= R2[0:7];
					R2[24:31] <= R3[0:7];
					R3[24:31] <= R4[0:7];
					R4[25:32] <= key;

					R1[0:22] <= R1[8:30];
					R2[0:23] <= R2[8:31];
					R3[0:23] <= R3[8:31];
					R4[0:24] <= R4[8:32];
				if (load_key) begin
					state <= State_Load_Key;
					end
				else if (load_iv)
					state <= State_Load_IV;
				else
					state <= State_Halt;
				end
			
			State_Load_IV: begin
				R1[23:30] <= {F1p1,F4p2,F3p3,F2p4,F1p5,F4p6,F3p7,F2p8};
				R2[24:31] <= {F2p1,F1p2,F4p3,F3p4,F2p5,F1p6,F4p7,F3p8};
				R3[24:31] <= {F3p1,F2p2,F1p3,F4p4,F3p5,F2p6,F1p7,F4p8};
				R4[25:32] <= {F4p1,F3p2,F2p3,F1p4,F4p5,F3p6,F2p7,F1p8};
				
				R1[0:22] <= R1[8:30];
				R2[0:23] <= R2[8:31];
				R3[0:23] <= R3[8:31];
				R4[0:24] <= R4[8:32];
				if (load_iv) begin
					state <= State_Load_IV;
					end
				else if (run)
					state <= State_Warm_Up;
				else
					state <= State_Halt;
				end
			
			State_Warm_Up: begin
				if (run) begin
					R1[23:30] <= {F1p1,F4p2,F3p3,F2p4,F1p5,F4p6,F3p7,F2p8};
					R2[24:31] <= {F2p1,F1p2,F4p3,F3p4,F2p5,F1p6,F4p7,F3p8};
					R3[24:31] <= {F3p1,F2p2,F1p3,F4p4,F3p5,F2p6,F1p7,F4p8};
					R4[25:32] <= {F4p1,F3p2,F2p3,F1p4,F4p5,F3p6,F2p7,F1p8};
					
					R1[0:22] <= R1[8:30];
					R2[0:23] <= R2[8:31];
					R3[0:23] <= R3[8:31];
					R4[0:24] <= R4[8:32];
					if (ready_counter < 3'b100) begin
						state <= State_Warm_Up;
						ready_counter <= ready_counter + 3'b01;
						end
					else if (ready_counter == 3'b100) begin
						warm_up_done <= 1'b1;
						state <= State_Gen_Output;
						end
					end
				else
					state <= State_Halt;
				end			
			
			State_Gen_Output:
				if (run) begin
					output_ready <= 1;
					stream_out <= R1[0:7]^R2[0:7]^R3[0:7]^R4[0:7];
					
					R1[23:30] <= {F1p1,F4p2,F3p3,F2p4,F1p5,F4p6,F3p7,F2p8};
					R2[24:31] <= {F2p1,F1p2,F4p3,F3p4,F2p5,F1p6,F4p7,F3p8};
					R3[24:31] <= {F3p1,F2p2,F1p3,F4p4,F3p5,F2p6,F1p7,F4p8};
					R4[25:32] <= {F4p1,F3p2,F2p3,F1p4,F4p5,F3p6,F2p7,F1p8};
					
					R1[0:22] <= R1[8:30];
					R2[0:23] <= R2[8:31];
					R3[0:23] <= R3[8:31];
					R4[0:24] <= R4[8:32];
					state <= State_Gen_Output;
					end
				else
					state <= State_Halt;
			
			State_Halt: 
				if (load_key)
					state <= State_Load_Key;
				else if (load_iv)
					state <= State_Load_IV;
				else if (run & ~warm_up_done)
					state <= State_Warm_Up;
				else if (run & warm_up_done)
					state <= State_Gen_Output;
				else
					state <= State_Halt;
				
			default state <= State_Halt;
			endcase


	//-----Feedback function of P1---------
	assign F1p1_ = R1[0] ^ R1[2] ^ R1[5] ^ R1[6] ^ R1[15] ^ R1[17] ^ R1[18] ^ R1[20] ^ R1[25] ^ (R1[8] & R1[18]) ^ (R1[8] & R1[20]) ^ (R1[12] & R1[21]) ^ (R1[14] & R1[19]) ^ (R1[17] & R1[21]) ^ ( R1[20] & R1[22]) ^ ( R1[4] & R1[12] & R1[22]) ^ ( R1[4] & R1[19] & R1[22]) ^ ( R1[7] & R1[20] & R1[21]) ^ ( R1[8] & R1[18] & R1[22]) ^ ( R1[8] & R1[20] & R1[22]) ^ ( R1[12] & R1[19] & R1[22]) ^ ( R1[20] & R1[21] & R1[22]) ^ ( R1[4] & R1[7] & R1[12] & R1[21]) ^ ( R1[4] & R1[7] & R1[19] & R1[21]) ^ ( R1[4] & R1[12] & R1[21] & R1[22]) ^ ( R1[4] & R1[19] & R1[21] & R1[22]) ^ ( R1[7] & R1[8] & R1[18] & R1[21]) ^ ( R1[7] & R1[8] & R1[20] & R1[21]) ^ ( R1[7] & R1[12] & R1[19] & R1[21]) ^ ( R1[8] & R1[18] & R1[21] & R1[22]) ^ ( R1[8] & R1[20] & R1[21] & R1[22]) ^ ( R1[12] & R1[19] & R1[21] & R1[22]);
	assign F2p1_ = R2[0] ^ R2[3] ^ R2[17] ^ R2[22] ^ R2[28]  ^ ( R2[2] & R2[13]) ^ ( R2[5] & R2[19]) ^ ( R2[7] & R2[19]) ^ ( R2[8] & R2[12]) ^ ( R2[8] & R2[13]) ^ ( R2[13] & R2[15]) ^ ( R2[2] & R2[12] & R2[13]) ^ ( R2[7] & R2[8] & R2[12]) ^ ( R2[7] & R2[8] & R2[14]) ^ ( R2[8] & R2[12] & R2[13]) ^ ( R2[2] & R2[7] & R2[12] & R2[13]) ^ ( R2[2] & R2[7] & R2[13] & R2[14]) ^ ( R2[4] & R2[11] & R2[12] & R2[24]) ^ ( R2[7] & R2[8] & R2[12] & R2[13]) ^ ( R2[7] & R2[8] & R2[13] & R2[14]) ^ ( R2[4] & R2[7] & R2[11] & R2[12] & R2[24]) ^ ( R2[4] & R2[7] & R2[11] & R2[14] & R2[24]);
	assign F3p1_ = R3[0] ^ R3[3] ^ R3[17] ^ R3[22] ^ R3[28]  ^ ( R3[2] & R3[13]) ^ ( R3[5] & R3[19]) ^ ( R3[7] & R3[19]) ^ ( R3[8] & R3[12]) ^ ( R3[8] & R3[13]) ^ ( R3[13] & R3[15]) ^ ( R3[2] & R3[12] & R3[13]) ^ ( R3[7] & R3[8] & R3[12]) ^ ( R3[7] & R3[8] & R3[14]) ^ ( R3[8] & R3[12] & R3[13]) ^ ( R3[2] & R3[7] & R3[12] & R3[13]) ^ ( R3[2] & R3[7] & R3[13] & R3[14]) ^ ( R3[4] & R3[11] & R3[12] & R3[24]) ^ ( R3[7] & R3[8] & R3[12] & R3[13]) ^ ( R3[7] & R3[8] & R3[13] & R3[14]) ^ ( R3[4] & R3[7] & R3[11] & R3[12] & R3[24]) ^ ( R3[4] & R3[7] & R3[11] & R3[14] & R3[24]);
	assign F4p1_ = R4[0] ^ R4[2] ^ R4[7] ^ R4[9] ^ R4[10] ^ R4[15] ^ R4[23] ^ R4[25] ^ R4[30] ^ ( R4[8] & R4[15]) ^ ( R4[12] & R4[16]) ^ ( R4[13] & R4[15]) ^ ( R4[13] & R4[25]) ^ ( R4[1] & R4[8] & R4[14]) ^ ( R4[1] & R4[8] & R4[18]) ^ ( R4[8] & R4[12] & R4[16]) ^ ( R4[8] & R4[14] & R4[18]) ^ ( R4[8] & R4[15] & R4[16]) ^ ( R4[8] & R4[15] & R4[17]) ^ ( R4[15] & R4[17] & R4[24]) ^ ( R4[1] & R4[8] & R4[14] & R4[17]) ^ ( R4[1] & R4[8] & R4[17] & R4[18]) ^ ( R4[1] & R4[14] & R4[17] & R4[24]) ^ ( R4[1] & R4[17] & R4[18] & R4[24]) ^ ( R4[8] & R4[12] & R4[16] & R4[17]) ^ ( R4[8] & R4[14] & R4[17] & R4[18]) ^ ( R4[8] & R4[15] & R4[16] & R4[17]) ^ ( R4[12] & R4[16] & R4[17] & R4[24]) ^ ( R4[14] & R4[17] & R4[18] & R4[24]) ^ ( R4[15] & R4[16] & R4[17] & R4[24]);
	
	assign F1p1 = (state == State_Load_IV)? F1p1_ ^ iv[0] : F1p1_;
	assign F2p1 = (state == State_Load_IV)? F2p1_ ^ iv[0] : F2p1_;
	assign F3p1 = (state == State_Load_IV)? F3p1_ ^ iv[0] : F3p1_;
	assign F4p1 = (state == State_Load_IV)? F4p1_ ^ iv[0] : F4p1_;

	//-----Feedback function of P2---------	
	assign F1p2_ = R1[0+1] ^ R1[2+1] ^ R1[5+1] ^ R1[6+1] ^ R1[15+1] ^ R1[17+1] ^ R1[18+1] ^ R1[20+1] ^ R1[25+1] ^ (R1[8+1] & R1[18+1]) ^ (R1[8+1] & R1[20+1]) ^ (R1[12+1] & R1[21+1]) ^ (R1[14+1] & R1[19+1]) ^ (R1[17+1] & R1[21+1]) ^ ( R1[20+1] & R1[22+1]) ^ ( R1[4+1] & R1[12+1] & R1[22+1]) ^ ( R1[4+1] & R1[19+1] & R1[22+1]) ^ ( R1[7+1] & R1[20+1] & R1[21+1]) ^ ( R1[8+1] & R1[18+1] & R1[22+1]) ^ ( R1[8+1] & R1[20+1] & R1[22+1]) ^ ( R1[12+1] & R1[19+1] & R1[22+1]) ^ ( R1[20+1] & R1[21+1] & R1[22+1]) ^ ( R1[4+1] & R1[7+1] & R1[12+1] & R1[21+1]) ^ ( R1[4+1] & R1[7+1] & R1[19+1] & R1[21+1]) ^ ( R1[4+1] & R1[12+1] & R1[21+1] & R1[22+1]) ^ ( R1[4+1] & R1[19+1] & R1[21+1] & R1[22+1]) ^ ( R1[7+1] & R1[8+1] & R1[18+1] & R1[21+1]) ^ ( R1[7+1] & R1[8+1] & R1[20+1] & R1[21+1]) ^ ( R1[7+1] & R1[12+1] & R1[19+1] & R1[21+1]) ^ ( R1[8+1] & R1[18+1] & R1[21+1] & R1[22+1]) ^ ( R1[8+1] & R1[20+1] & R1[21+1] & R1[22+1]) ^ ( R1[12+1] & R1[19+1] & R1[21+1] & R1[22+1]);
	assign F2p2_ = R2[0+1] ^ R2[3+1] ^ R2[17+1] ^ R2[22+1] ^ R2[28+1]  ^ ( R2[2+1] & R2[13+1]) ^ ( R2[5+1] & R2[19+1]) ^ ( R2[7+1] & R2[19+1]) ^ ( R2[8+1] & R2[12+1]) ^ ( R2[8+1] & R2[13+1]) ^ ( R2[13+1] & R2[15+1]) ^ ( R2[2+1] & R2[12+1] & R2[13+1]) ^ ( R2[7+1] & R2[8+1] & R2[12+1]) ^ ( R2[7+1] & R2[8+1] & R2[14+1]) ^ ( R2[8+1] & R2[12+1] & R2[13+1]) ^ ( R2[2+1] & R2[7+1] & R2[12+1] & R2[13+1]) ^ ( R2[2+1] & R2[7+1] & R2[13+1] & R2[14+1]) ^ ( R2[4+1] & R2[11+1] & R2[12+1] & R2[24+1]) ^ ( R2[7+1] & R2[8+1] & R2[12+1] & R2[13+1]) ^ ( R2[7+1] & R2[8+1] & R2[13+1] & R2[14+1]) ^ ( R2[4+1] & R2[7+1] & R2[11+1] & R2[12+1] & R2[24+1]) ^ ( R2[4+1] & R2[7+1] & R2[11+1] & R2[14+1] & R2[24+1]);
	assign F3p2_ = R3[0+1] ^ R3[3+1] ^ R3[17+1] ^ R3[22+1] ^ R3[28+1]  ^ ( R3[2+1] & R3[13+1]) ^ ( R3[5+1] & R3[19+1]) ^ ( R3[7+1] & R3[19+1]) ^ ( R3[8+1] & R3[12+1]) ^ ( R3[8+1] & R3[13+1]) ^ ( R3[13+1] & R3[15+1]) ^ ( R3[2+1] & R3[12+1] & R3[13+1]) ^ ( R3[7+1] & R3[8+1] & R3[12+1]) ^ ( R3[7+1] & R3[8+1] & R3[14+1]) ^ ( R3[8+1] & R3[12+1] & R3[13+1]) ^ ( R3[2+1] & R3[7+1] & R3[12+1] & R3[13+1]) ^ ( R3[2+1] & R3[7+1] & R3[13+1] & R3[14+1]) ^ ( R3[4+1] & R3[11+1] & R3[12+1] & R3[24+1]) ^ ( R3[7+1] & R3[8+1] & R3[12+1] & R3[13+1]) ^ ( R3[7+1] & R3[8+1] & R3[13+1] & R3[14+1]) ^ ( R3[4+1] & R3[7+1] & R3[11+1] & R3[12+1] & R3[24+1]) ^ ( R3[4+1] & R3[7+1] & R3[11+1] & R3[14+1] & R3[24+1]);
	assign F4p2_ = R4[0+1] ^ R4[2+1] ^ R4[7+1] ^ R4[9+1] ^ R4[10+1] ^ R4[15+1] ^ R4[23+1] ^ R4[25+1] ^ R4[30+1] ^ ( R4[8+1] & R4[15+1]) ^ ( R4[12+1] & R4[16+1]) ^ ( R4[13+1] & R4[15+1]) ^ ( R4[13+1] & R4[25+1]) ^ ( R4[1+1] & R4[8+1] & R4[14+1]) ^ ( R4[1+1] & R4[8+1] & R4[18+1]) ^ ( R4[8+1] & R4[12+1] & R4[16+1]) ^ ( R4[8+1] & R4[14+1] & R4[18+1]) ^ ( R4[8+1] & R4[15+1] & R4[16+1]) ^ ( R4[8+1] & R4[15+1] & R4[17+1]) ^ ( R4[15+1] & R4[17+1] & R4[24+1]) ^ ( R4[1+1] & R4[8+1] & R4[14+1] & R4[17+1]) ^ ( R4[1+1] & R4[8+1] & R4[17+1] & R4[18+1]) ^ ( R4[1+1] & R4[14+1] & R4[17+1] & R4[24+1]) ^ ( R4[1+1] & R4[17+1] & R4[18+1] & R4[24+1]) ^ ( R4[8+1] & R4[12+1] & R4[16+1] & R4[17+1]) ^ ( R4[8+1] & R4[14+1] & R4[17+1] & R4[18+1]) ^ ( R4[8+1] & R4[15+1] & R4[16+1] & R4[17+1]) ^ ( R4[12+1] & R4[16+1] & R4[17+1] & R4[24+1]) ^ ( R4[14+1] & R4[17+1] & R4[18+1] & R4[24+1]) ^ ( R4[15+1] & R4[16+1] & R4[17+1] & R4[24+1]);
	
	assign F1p2 = (state == State_Load_IV)? F1p2_ ^ iv[0+1] : F1p2_;
	assign F2p2 = (state == State_Load_IV)? F2p2_ ^ iv[0+1] : F2p2_;
	assign F3p2 = (state == State_Load_IV)? F3p2_ ^ iv[0+1] : F3p2_;
	assign F4p2 = (state == State_Load_IV)? F4p2_ ^ iv[0+1] : F4p2_;
	
	//-----Feedback function of P3---------	
	assign F1p3_ = R1[0+2] ^ R1[2+2] ^ R1[5+2] ^ R1[6+2] ^ R1[15+2] ^ R1[17+2] ^ R1[18+2] ^ R1[20+2] ^ R1[25+2] ^ (R1[8+2] & R1[18+2]) ^ (R1[8+2] & R1[20+2]) ^ (R1[12+2] & R1[21+2]) ^ (R1[14+2] & R1[19+2]) ^ (R1[17+2] & R1[21+2]) ^ ( R1[20+2] & R1[22+2]) ^ ( R1[4+2] & R1[12+2] & R1[22+2]) ^ ( R1[4+2] & R1[19+2] & R1[22+2]) ^ ( R1[7+2] & R1[20+2] & R1[21+2]) ^ ( R1[8+2] & R1[18+2] & R1[22+2]) ^ ( R1[8+2] & R1[20+2] & R1[22+2]) ^ ( R1[12+2] & R1[19+2] & R1[22+2]) ^ ( R1[20+2] & R1[21+2] & R1[22+2]) ^ ( R1[4+2] & R1[7+2] & R1[12+2] & R1[21+2]) ^ ( R1[4+2] & R1[7+2] & R1[19+2] & R1[21+2]) ^ ( R1[4+2] & R1[12+2] & R1[21+2] & R1[22+2]) ^ ( R1[4+2] & R1[19+2] & R1[21+2] & R1[22+2]) ^ ( R1[7+2] & R1[8+2] & R1[18+2] & R1[21+2]) ^ ( R1[7+2] & R1[8+2] & R1[20+2] & R1[21+2]) ^ ( R1[7+2] & R1[12+2] & R1[19+2] & R1[21+2]) ^ ( R1[8+2] & R1[18+2] & R1[21+2] & R1[22+2]) ^ ( R1[8+2] & R1[20+2] & R1[21+2] & R1[22+2]) ^ ( R1[12+2] & R1[19+2] & R1[21+2] & R1[22+2]);
	assign F2p3_ = R2[0+2] ^ R2[3+2] ^ R2[17+2] ^ R2[22+2] ^ R2[28+2]  ^ ( R2[2+2] & R2[13+2]) ^ ( R2[5+2] & R2[19+2]) ^ ( R2[7+2] & R2[19+2]) ^ ( R2[8+2] & R2[12+2]) ^ ( R2[8+2] & R2[13+2]) ^ ( R2[13+2] & R2[15+2]) ^ ( R2[2+2] & R2[12+2] & R2[13+2]) ^ ( R2[7+2] & R2[8+2] & R2[12+2]) ^ ( R2[7+2] & R2[8+2] & R2[14+2]) ^ ( R2[8+2] & R2[12+2] & R2[13+2]) ^ ( R2[2+2] & R2[7+2] & R2[12+2] & R2[13+2]) ^ ( R2[2+2] & R2[7+2] & R2[13+2] & R2[14+2]) ^ ( R2[4+2] & R2[11+2] & R2[12+2] & R2[24+2]) ^ ( R2[7+2] & R2[8+2] & R2[12+2] & R2[13+2]) ^ ( R2[7+2] & R2[8+2] & R2[13+2] & R2[14+2]) ^ ( R2[4+2] & R2[7+2] & R2[11+2] & R2[12+2] & R2[24+2]) ^ ( R2[4+2] & R2[7+2] & R2[11+2] & R2[14+2] & R2[24+2]);
	assign F3p3_ = R3[0+2] ^ R3[3+2] ^ R3[17+2] ^ R3[22+2] ^ R3[28+2]  ^ ( R3[2+2] & R3[13+2]) ^ ( R3[5+2] & R3[19+2]) ^ ( R3[7+2] & R3[19+2]) ^ ( R3[8+2] & R3[12+2]) ^ ( R3[8+2] & R3[13+2]) ^ ( R3[13+2] & R3[15+2]) ^ ( R3[2+2] & R3[12+2] & R3[13+2]) ^ ( R3[7+2] & R3[8+2] & R3[12+2]) ^ ( R3[7+2] & R3[8+2] & R3[14+2]) ^ ( R3[8+2] & R3[12+2] & R3[13+2]) ^ ( R3[2+2] & R3[7+2] & R3[12+2] & R3[13+2]) ^ ( R3[2+2] & R3[7+2] & R3[13+2] & R3[14+2]) ^ ( R3[4+2] & R3[11+2] & R3[12+2] & R3[24+2]) ^ ( R3[7+2] & R3[8+2] & R3[12+2] & R3[13+2]) ^ ( R3[7+2] & R3[8+2] & R3[13+2] & R3[14+2]) ^ ( R3[4+2] & R3[7+2] & R3[11+2] & R3[12+2] & R3[24+2]) ^ ( R3[4+2] & R3[7+2] & R3[11+2] & R3[14+2] & R3[24+2]);
	assign F4p3_ = R4[0+2] ^ R4[2+2] ^ R4[7+2] ^ R4[9+2] ^ R4[10+2] ^ R4[15+2] ^ R4[23+2] ^ R4[25+2] ^ R4[30+2] ^ ( R4[8+2] & R4[15+2]) ^ ( R4[12+2] & R4[16+2]) ^ ( R4[13+2] & R4[15+2]) ^ ( R4[13+2] & R4[25+2]) ^ ( R4[1+2] & R4[8+2] & R4[14+2]) ^ ( R4[1+2] & R4[8+2] & R4[18+2]) ^ ( R4[8+2] & R4[12+2] & R4[16+2]) ^ ( R4[8+2] & R4[14+2] & R4[18+2]) ^ ( R4[8+2] & R4[15+2] & R4[16+2]) ^ ( R4[8+2] & R4[15+2] & R4[17+2]) ^ ( R4[15+2] & R4[17+2] & R4[24+2]) ^ ( R4[1+2] & R4[8+2] & R4[14+2] & R4[17+2]) ^ ( R4[1+2] & R4[8+2] & R4[17+2] & R4[18+2]) ^ ( R4[1+2] & R4[14+2] & R4[17+2] & R4[24+2]) ^ ( R4[1+2] & R4[17+2] & R4[18+2] & R4[24+2]) ^ ( R4[8+2] & R4[12+2] & R4[16+2] & R4[17+2]) ^ ( R4[8+2] & R4[14+2] & R4[17+2] & R4[18+2]) ^ ( R4[8+2] & R4[15+2] & R4[16+2] & R4[17+2]) ^ ( R4[12+2] & R4[16+2] & R4[17+2] & R4[24+2]) ^ ( R4[14+2] & R4[17+2] & R4[18+2] & R4[24+2]) ^ ( R4[15+2] & R4[16+2] & R4[17+2] & R4[24+2]);
	
	assign F1p3 = (state == State_Load_IV)? F1p3_ ^ iv[0+2] : F1p3_;
	assign F2p3 = (state == State_Load_IV)? F2p3_ ^ iv[0+2] : F2p3_;
	assign F3p3 = (state == State_Load_IV)? F3p3_ ^ iv[0+2] : F3p3_;
	assign F4p3 = (state == State_Load_IV)? F4p3_ ^ iv[0+2] : F4p3_;	
	
		//-----Feedback function of P4---------	
	assign F1p4_ = R1[0+3] ^ R1[2+3] ^ R1[5+3] ^ R1[6+3] ^ R1[15+3] ^ R1[17+3] ^ R1[18+3] ^ R1[20+3] ^ R1[25+3] ^ (R1[8+3] & R1[18+3]) ^ (R1[8+3] & R1[20+3]) ^ (R1[12+3] & R1[21+3]) ^ (R1[14+3] & R1[19+3]) ^ (R1[17+3] & R1[21+3]) ^ ( R1[20+3] & R1[22+3]) ^ ( R1[4+3] & R1[12+3] & R1[22+3]) ^ ( R1[4+3] & R1[19+3] & R1[22+3]) ^ ( R1[7+3] & R1[20+3] & R1[21+3]) ^ ( R1[8+3] & R1[18+3] & R1[22+3]) ^ ( R1[8+3] & R1[20+3] & R1[22+3]) ^ ( R1[12+3] & R1[19+3] & R1[22+3]) ^ ( R1[20+3] & R1[21+3] & R1[22+3]) ^ ( R1[4+3] & R1[7+3] & R1[12+3] & R1[21+3]) ^ ( R1[4+3] & R1[7+3] & R1[19+3] & R1[21+3]) ^ ( R1[4+3] & R1[12+3] & R1[21+3] & R1[22+3]) ^ ( R1[4+3] & R1[19+3] & R1[21+3] & R1[22+3]) ^ ( R1[7+3] & R1[8+3] & R1[18+3] & R1[21+3]) ^ ( R1[7+3] & R1[8+3] & R1[20+3] & R1[21+3]) ^ ( R1[7+3] & R1[12+3] & R1[19+3] & R1[21+3]) ^ ( R1[8+3] & R1[18+3] & R1[21+3] & R1[22+3]) ^ ( R1[8+3] & R1[20+3] & R1[21+3] & R1[22+3]) ^ ( R1[12+3] & R1[19+3] & R1[21+3] & R1[22+3]);
	assign F2p4_ = R2[0+3] ^ R2[3+3] ^ R2[17+3] ^ R2[22+3] ^ R2[28+3]  ^ ( R2[2+3] & R2[13+3]) ^ ( R2[5+3] & R2[19+3]) ^ ( R2[7+3] & R2[19+3]) ^ ( R2[8+3] & R2[12+3]) ^ ( R2[8+3] & R2[13+3]) ^ ( R2[13+3] & R2[15+3]) ^ ( R2[2+3] & R2[12+3] & R2[13+3]) ^ ( R2[7+3] & R2[8+3] & R2[12+3]) ^ ( R2[7+3] & R2[8+3] & R2[14+3]) ^ ( R2[8+3] & R2[12+3] & R2[13+3]) ^ ( R2[2+3] & R2[7+3] & R2[12+3] & R2[13+3]) ^ ( R2[2+3] & R2[7+3] & R2[13+3] & R2[14+3]) ^ ( R2[4+3] & R2[11+3] & R2[12+3] & R2[24+3]) ^ ( R2[7+3] & R2[8+3] & R2[12+3] & R2[13+3]) ^ ( R2[7+3] & R2[8+3] & R2[13+3] & R2[14+3]) ^ ( R2[4+3] & R2[7+3] & R2[11+3] & R2[12+3] & R2[24+3]) ^ ( R2[4+3] & R2[7+3] & R2[11+3] & R2[14+3] & R2[24+3]);
	assign F3p4_ = R3[0+3] ^ R3[3+3] ^ R3[17+3] ^ R3[22+3] ^ R3[28+3]  ^ ( R3[2+3] & R3[13+3]) ^ ( R3[5+3] & R3[19+3]) ^ ( R3[7+3] & R3[19+3]) ^ ( R3[8+3] & R3[12+3]) ^ ( R3[8+3] & R3[13+3]) ^ ( R3[13+3] & R3[15+3]) ^ ( R3[2+3] & R3[12+3] & R3[13+3]) ^ ( R3[7+3] & R3[8+3] & R3[12+3]) ^ ( R3[7+3] & R3[8+3] & R3[14+3]) ^ ( R3[8+3] & R3[12+3] & R3[13+3]) ^ ( R3[2+3] & R3[7+3] & R3[12+3] & R3[13+3]) ^ ( R3[2+3] & R3[7+3] & R3[13+3] & R3[14+3]) ^ ( R3[4+3] & R3[11+3] & R3[12+3] & R3[24+3]) ^ ( R3[7+3] & R3[8+3] & R3[12+3] & R3[13+3]) ^ ( R3[7+3] & R3[8+3] & R3[13+3] & R3[14+3]) ^ ( R3[4+3] & R3[7+3] & R3[11+3] & R3[12+3] & R3[24+3]) ^ ( R3[4+3] & R3[7+3] & R3[11+3] & R3[14+3] & R3[24+3]);
	assign F4p4_ = R4[0+3] ^ R4[2+3] ^ R4[7+3] ^ R4[9+3] ^ R4[10+3] ^ R4[15+3] ^ R4[23+3] ^ R4[25+3] ^ F4p1 ^ ( R4[8+3] & R4[15+3]) ^ ( R4[12+3] & R4[16+3]) ^ ( R4[13+3] & R4[15+3]) ^ ( R4[13+3] & R4[25+3]) ^ ( R4[1+3] & R4[8+3] & R4[14+3]) ^ ( R4[1+3] & R4[8+3] & R4[18+3]) ^ ( R4[8+3] & R4[12+3] & R4[16+3]) ^ ( R4[8+3] & R4[14+3] & R4[18+3]) ^ ( R4[8+3] & R4[15+3] & R4[16+3]) ^ ( R4[8+3] & R4[15+3] & R4[17+3]) ^ ( R4[15+3] & R4[17+3] & R4[24+3]) ^ ( R4[1+3] & R4[8+3] & R4[14+3] & R4[17+3]) ^ ( R4[1+3] & R4[8+3] & R4[17+3] & R4[18+3]) ^ ( R4[1+3] & R4[14+3] & R4[17+3] & R4[24+3]) ^ ( R4[1+3] & R4[17+3] & R4[18+3] & R4[24+3]) ^ ( R4[8+3] & R4[12+3] & R4[16+3] & R4[17+3]) ^ ( R4[8+3] & R4[14+3] & R4[17+3] & R4[18+3]) ^ ( R4[8+3] & R4[15+3] & R4[16+3] & R4[17+3]) ^ ( R4[12+3] & R4[16+3] & R4[17+3] & R4[24+3]) ^ ( R4[14+3] & R4[17+3] & R4[18+3] & R4[24+3]) ^ ( R4[15+3] & R4[16+3] & R4[17+3] & R4[24+3]);
	
	assign F1p4 = (state == State_Load_IV)? F1p4_ ^ iv[0+3] : F1p4_;
	assign F2p4 = (state == State_Load_IV)? F2p4_ ^ iv[0+3] : F2p4_;
	assign F3p4 = (state == State_Load_IV)? F3p4_ ^ iv[0+3] : F3p4_;
	assign F4p4 = (state == State_Load_IV)? F4p4_ ^ iv[0+3] : F4p4_;	

	//-----Feedback function of P5---------
	assign F1p5_ = R1[0+4] ^ R1[2+4] ^ R1[5+4] ^ R1[6+4] ^ R1[15+4] ^ R1[17+4] ^ R1[18+4] ^ R1[20+4] ^ R1[25+4] ^ (R1[8+4] & R1[18+4]) ^ (R1[8+4] & R1[20+4]) ^ (R1[12+4] & R1[21+4]) ^ (R1[14+4] & R1[19+4]) ^ (R1[17+4] & R1[21+4]) ^ ( R1[20+4] & R1[22+4]) ^ ( R1[4+4] & R1[12+4] & R1[22+4]) ^ ( R1[4+4] & R1[19+4] & R1[22+4]) ^ ( R1[7+4] & R1[20+4] & R1[21+4]) ^ ( R1[8+4] & R1[18+4] & R1[22+4]) ^ ( R1[8+4] & R1[20+4] & R1[22+4]) ^ ( R1[12+4] & R1[19+4] & R1[22+4]) ^ ( R1[20+4] & R1[21+4] & R1[22+4]) ^ ( R1[4+4] & R1[7+4] & R1[12+4] & R1[21+4]) ^ ( R1[4+4] & R1[7+4] & R1[19+4] & R1[21+4]) ^ ( R1[4+4] & R1[12+4] & R1[21+4] & R1[22+4]) ^ ( R1[4+4] & R1[19+4] & R1[21+4] & R1[22+4]) ^ ( R1[7+4] & R1[8+4] & R1[18+4] & R1[21+4]) ^ ( R1[7+4] & R1[8+4] & R1[20+4] & R1[21+4]) ^ ( R1[7+4] & R1[12+4] & R1[19+4] & R1[21+4]) ^ ( R1[8+4] & R1[18+4] & R1[21+4] & R1[22+4]) ^ ( R1[8+4] & R1[20+4] & R1[21+4] & R1[22+4]) ^ ( R1[12+4] & R1[19+4] & R1[21+4] & R1[22+4]);
	assign F2p5_ = R2[0+4] ^ R2[3+4] ^ R2[17+4] ^ R2[22+4] ^ F2p1  ^ ( R2[2+4] & R2[13+4]) ^ ( R2[5+4] & R2[19+4]) ^ ( R2[7+4] & R2[19+4]) ^ ( R2[8+4] & R2[12+4]) ^ ( R2[8+4] & R2[13+4]) ^ ( R2[13+4] & R2[15+4]) ^ ( R2[2+4] & R2[12+4] & R2[13+4]) ^ ( R2[7+4] & R2[8+4] & R2[12+4]) ^ ( R2[7+4] & R2[8+4] & R2[14+4]) ^ ( R2[8+4] & R2[12+4] & R2[13+4]) ^ ( R2[2+4] & R2[7+4] & R2[12+4] & R2[13+4]) ^ ( R2[2+4] & R2[7+4] & R2[13+4] & R2[14+4]) ^ ( R2[4+4] & R2[11+4] & R2[12+4] & R2[24+4]) ^ ( R2[7+4] & R2[8+4] & R2[12+4] & R2[13+4]) ^ ( R2[7+4] & R2[8+4] & R2[13+4] & R2[14+4]) ^ ( R2[4+4] & R2[7+4] & R2[11+4] & R2[12+4] & R2[24+4]) ^ ( R2[4+4] & R2[7+4] & R2[11+4] & R2[14+4] & R2[24+4]);
	assign F3p5_ = R3[0+4] ^ R3[3+4] ^ R3[17+4] ^ R3[22+4] ^ F3p1  ^ ( R3[2+4] & R3[13+4]) ^ ( R3[5+4] & R3[19+4]) ^ ( R3[7+4] & R3[19+4]) ^ ( R3[8+4] & R3[12+4]) ^ ( R3[8+4] & R3[13+4]) ^ ( R3[13+4] & R3[15+4]) ^ ( R3[2+4] & R3[12+4] & R3[13+4]) ^ ( R3[7+4] & R3[8+4] & R3[12+4]) ^ ( R3[7+4] & R3[8+4] & R3[14+4]) ^ ( R3[8+4] & R3[12+4] & R3[13+4]) ^ ( R3[2+4] & R3[7+4] & R3[12+4] & R3[13+4]) ^ ( R3[2+4] & R3[7+4] & R3[13+4] & R3[14+4]) ^ ( R3[4+4] & R3[11+4] & R3[12+4] & R3[24+4]) ^ ( R3[7+4] & R3[8+4] & R3[12+4] & R3[13+4]) ^ ( R3[7+4] & R3[8+4] & R3[13+4] & R3[14+4]) ^ ( R3[4+4] & R3[7+4] & R3[11+4] & R3[12+4] & R3[24+4]) ^ ( R3[4+4] & R3[7+4] & R3[11+4] & R3[14+4] & R3[24+4]);
	assign F4p5_ = R4[0+4] ^ R4[2+4] ^ R4[7+4] ^ R4[9+4] ^ R4[10+4] ^ R4[15+4] ^ R4[23+4] ^ R4[25+4] ^ F3p2 ^ ( R4[8+4] & R4[15+4]) ^ ( R4[12+4] & R4[16+4]) ^ ( R4[13+4] & R4[15+4]) ^ ( R4[13+4] & R4[25+4]) ^ ( R4[1+4] & R4[8+4] & R4[14+4]) ^ ( R4[1+4] & R4[8+4] & R4[18+4]) ^ ( R4[8+4] & R4[12+4] & R4[16+4]) ^ ( R4[8+4] & R4[14+4] & R4[18+4]) ^ ( R4[8+4] & R4[15+4] & R4[16+4]) ^ ( R4[8+4] & R4[15+4] & R4[17+4]) ^ ( R4[15+4] & R4[17+4] & R4[24+4]) ^ ( R4[1+4] & R4[8+4] & R4[14+4] & R4[17+4]) ^ ( R4[1+4] & R4[8+4] & R4[17+4] & R4[18+4]) ^ ( R4[1+4] & R4[14+4] & R4[17+4] & R4[24+4]) ^ ( R4[1+4] & R4[17+4] & R4[18+4] & R4[24+4]) ^ ( R4[8+4] & R4[12+4] & R4[16+4] & R4[17+4]) ^ ( R4[8+4] & R4[14+4] & R4[17+4] & R4[18+4]) ^ ( R4[8+4] & R4[15+4] & R4[16+4] & R4[17+4]) ^ ( R4[12+4] & R4[16+4] & R4[17+4] & R4[24+4]) ^ ( R4[14+4] & R4[17+4] & R4[18+4] & R4[24+4]) ^ ( R4[15+4] & R4[16+4] & R4[17+4] & R4[24+4]);
	
	assign F1p5 = (state == State_Load_IV)? F1p5_ ^ iv[0+4] : F1p5_;
	assign F2p5 = (state == State_Load_IV)? F2p5_ ^ iv[0+4] : F2p5_;
	assign F3p5 = (state == State_Load_IV)? F3p5_ ^ iv[0+4] : F3p5_;
	assign F4p5 = (state == State_Load_IV)? F4p5_ ^ iv[0+4] : F4p5_;
	
	//-----Feedback function of P6---------
	assign F1p6_ = R1[0+5] ^ R1[2+5] ^ R1[5+5] ^ R1[6+5] ^ R1[15+5] ^ R1[17+5] ^ R1[18+5] ^ R1[20+5] ^ R1[25+5] ^ (R1[8+5] & R1[18+5]) ^ (R1[8+5] & R1[20+5]) ^ (R1[12+5] & R1[21+5]) ^ (R1[14+5] & R1[19+5]) ^ (R1[17+5] & R1[21+5]) ^ ( R1[20+5] & R1[22+5]) ^ ( R1[4+5] & R1[12+5] & R1[22+5]) ^ ( R1[4+5] & R1[19+5] & R1[22+5]) ^ ( R1[7+5] & R1[20+5] & R1[21+5]) ^ ( R1[8+5] & R1[18+5] & R1[22+5]) ^ ( R1[8+5] & R1[20+5] & R1[22+5]) ^ ( R1[12+5] & R1[19+5] & R1[22+5]) ^ ( R1[20+5] & R1[21+5] & R1[22+5]) ^ ( R1[4+5] & R1[7+5] & R1[12+5] & R1[21+5]) ^ ( R1[4+5] & R1[7+5] & R1[19+5] & R1[21+5]) ^ ( R1[4+5] & R1[12+5] & R1[21+5] & R1[22+5]) ^ ( R1[4+5] & R1[19+5] & R1[21+5] & R1[22+5]) ^ ( R1[7+5] & R1[8+5] & R1[18+5] & R1[21+5]) ^ ( R1[7+5] & R1[8+5] & R1[20+5] & R1[21+5]) ^ ( R1[7+5] & R1[12+5] & R1[19+5] & R1[21+5]) ^ ( R1[8+5] & R1[18+5] & R1[21+5] & R1[22+5]) ^ ( R1[8+5] & R1[20+5] & R1[21+5] & R1[22+5]) ^ ( R1[12+5] & R1[19+5] & R1[21+5] & R1[22+5]);
	assign F2p6_ = R2[0+5] ^ R2[3+5] ^ R2[17+5] ^ R2[22+5] ^ F1p2  ^ ( R2[2+5] & R2[13+5]) ^ ( R2[5+5] & R2[19+5]) ^ ( R2[7+5] & R2[19+5]) ^ ( R2[8+5] & R2[12+5]) ^ ( R2[8+5] & R2[13+5]) ^ ( R2[13+5] & R2[15+5]) ^ ( R2[2+5] & R2[12+5] & R2[13+5]) ^ ( R2[7+5] & R2[8+5] & R2[12+5]) ^ ( R2[7+5] & R2[8+5] & R2[14+5]) ^ ( R2[8+5] & R2[12+5] & R2[13+5]) ^ ( R2[2+5] & R2[7+5] & R2[12+5] & R2[13+5]) ^ ( R2[2+5] & R2[7+5] & R2[13+5] & R2[14+5]) ^ ( R2[4+5] & R2[11+5] & R2[12+5] & R2[24+5]) ^ ( R2[7+5] & R2[8+5] & R2[12+5] & R2[13+5]) ^ ( R2[7+5] & R2[8+5] & R2[13+5] & R2[14+5]) ^ ( R2[4+5] & R2[7+5] & R2[11+5] & R2[12+5] & R2[24+5]) ^ ( R2[4+5] & R2[7+5] & R2[11+5] & R2[14+5] & R2[24+5]);
	assign F3p6_ = R3[0+5] ^ R3[3+5] ^ R3[17+5] ^ R3[22+5] ^ F2p2  ^ ( R3[2+5] & R3[13+5]) ^ ( R3[5+5] & R3[19+5]) ^ ( R3[7+5] & R3[19+5]) ^ ( R3[8+5] & R3[12+5]) ^ ( R3[8+5] & R3[13+5]) ^ ( R3[13+5] & R3[15+5]) ^ ( R3[2+5] & R3[12+5] & R3[13+5]) ^ ( R3[7+5] & R3[8+5] & R3[12+5]) ^ ( R3[7+5] & R3[8+5] & R3[14+5]) ^ ( R3[8+5] & R3[12+5] & R3[13+5]) ^ ( R3[2+5] & R3[7+5] & R3[12+5] & R3[13+5]) ^ ( R3[2+5] & R3[7+5] & R3[13+5] & R3[14+5]) ^ ( R3[4+5] & R3[11+5] & R3[12+5] & R3[24+5]) ^ ( R3[7+5] & R3[8+5] & R3[12+5] & R3[13+5]) ^ ( R3[7+5] & R3[8+5] & R3[13+5] & R3[14+5]) ^ ( R3[4+5] & R3[7+5] & R3[11+5] & R3[12+5] & R3[24+5]) ^ ( R3[4+5] & R3[7+5] & R3[11+5] & R3[14+5] & R3[24+5]);
	assign F4p6_ = R4[0+5] ^ R4[2+5] ^ R4[7+5] ^ R4[9+5] ^ R4[10+5] ^ R4[15+5] ^ R4[23+5] ^ R4[25+5] ^ F2p3 ^ ( R4[8+5] & R4[15+5]) ^ ( R4[12+5] & R4[16+5]) ^ ( R4[13+5] & R4[15+5]) ^ ( R4[13+5] & R4[25+5]) ^ ( R4[1+5] & R4[8+5] & R4[14+5]) ^ ( R4[1+5] & R4[8+5] & R4[18+5]) ^ ( R4[8+5] & R4[12+5] & R4[16+5]) ^ ( R4[8+5] & R4[14+5] & R4[18+5]) ^ ( R4[8+5] & R4[15+5] & R4[16+5]) ^ ( R4[8+5] & R4[15+5] & R4[17+5]) ^ ( R4[15+5] & R4[17+5] & R4[24+5]) ^ ( R4[1+5] & R4[8+5] & R4[14+5] & R4[17+5]) ^ ( R4[1+5] & R4[8+5] & R4[17+5] & R4[18+5]) ^ ( R4[1+5] & R4[14+5] & R4[17+5] & R4[24+5]) ^ ( R4[1+5] & R4[17+5] & R4[18+5] & R4[24+5]) ^ ( R4[8+5] & R4[12+5] & R4[16+5] & R4[17+5]) ^ ( R4[8+5] & R4[14+5] & R4[17+5] & R4[18+5]) ^ ( R4[8+5] & R4[15+5] & R4[16+5] & R4[17+5]) ^ ( R4[12+5] & R4[16+5] & R4[17+5] & R4[24+5]) ^ ( R4[14+5] & R4[17+5] & R4[18+5] & R4[24+5]) ^ ( R4[15+5] & R4[16+5] & R4[17+5] & R4[24+5]);

	assign F1p6 = (state == State_Load_IV)? F1p6_ ^ iv[0+5] : F1p6_;
	assign F2p6 = (state == State_Load_IV)? F2p6_ ^ iv[0+5] : F2p6_;
	assign F3p6 = (state == State_Load_IV)? F3p6_ ^ iv[0+5] : F3p6_;
	assign F4p6 = (state == State_Load_IV)? F4p6_ ^ iv[0+5] : F4p6_;
	
	//-----Feedback function of P7---------
	assign F1p7_ = R1[0+6] ^ R1[2+6] ^ R1[5+6] ^ R1[6+6] ^ R1[15+6] ^ R1[17+6] ^ R1[18+6] ^ R1[20+6] ^ F1p1 ^ (R1[8+6] & R1[18+6]) ^ (R1[8+6] & R1[20+6]) ^ (R1[12+6] & R1[21+6]) ^ (R1[14+6] & R1[19+6]) ^ (R1[17+6] & R1[21+6]) ^ ( R1[20+6] & R1[22+6]) ^ ( R1[4+6] & R1[12+6] & R1[22+6]) ^ ( R1[4+6] & R1[19+6] & R1[22+6]) ^ ( R1[7+6] & R1[20+6] & R1[21+6]) ^ ( R1[8+6] & R1[18+6] & R1[22+6]) ^ ( R1[8+6] & R1[20+6] & R1[22+6]) ^ ( R1[12+6] & R1[19+6] & R1[22+6]) ^ ( R1[20+6] & R1[21+6] & R1[22+6]) ^ ( R1[4+6] & R1[7+6] & R1[12+6] & R1[21+6]) ^ ( R1[4+6] & R1[7+6] & R1[19+6] & R1[21+6]) ^ ( R1[4+6] & R1[12+6] & R1[21+6] & R1[22+6]) ^ ( R1[4+6] & R1[19+6] & R1[21+6] & R1[22+6]) ^ ( R1[7+6] & R1[8+6] & R1[18+6] & R1[21+6]) ^ ( R1[7+6] & R1[8+6] & R1[20+6] & R1[21+6]) ^ ( R1[7+6] & R1[12+6] & R1[19+6] & R1[21+6]) ^ ( R1[8+6] & R1[18+6] & R1[21+6] & R1[22+6]) ^ ( R1[8+6] & R1[20+6] & R1[21+6] & R1[22+6]) ^ ( R1[12+6] & R1[19+6] & R1[21+6] & R1[22+6]);
	assign F2p7_ = R2[0+6] ^ R2[3+6] ^ R2[17+6] ^ R2[22+6] ^ F4p3  ^ ( R2[2+6] & R2[13+6]) ^ ( R2[5+6] & R2[19+6]) ^ ( R2[7+6] & R2[19+6]) ^ ( R2[8+6] & R2[12+6]) ^ ( R2[8+6] & R2[13+6]) ^ ( R2[13+6] & R2[15+6]) ^ ( R2[2+6] & R2[12+6] & R2[13+6]) ^ ( R2[7+6] & R2[8+6] & R2[12+6]) ^ ( R2[7+6] & R2[8+6] & R2[14+6]) ^ ( R2[8+6] & R2[12+6] & R2[13+6]) ^ ( R2[2+6] & R2[7+6] & R2[12+6] & R2[13+6]) ^ ( R2[2+6] & R2[7+6] & R2[13+6] & R2[14+6]) ^ ( R2[4+6] & R2[11+6] & R2[12+6] & R2[24+6]) ^ ( R2[7+6] & R2[8+6] & R2[12+6] & R2[13+6]) ^ ( R2[7+6] & R2[8+6] & R2[13+6] & R2[14+6]) ^ ( R2[4+6] & R2[7+6] & R2[11+6] & R2[12+6] & R2[24+6]) ^ ( R2[4+6] & R2[7+6] & R2[11+6] & R2[14+6] & R2[24+6]);
	assign F3p7_ = R3[0+6] ^ R3[3+6] ^ R3[17+6] ^ R3[22+6] ^ F1p3  ^ ( R3[2+6] & R3[13+6]) ^ ( R3[5+6] & R3[19+6]) ^ ( R3[7+6] & R3[19+6]) ^ ( R3[8+6] & R3[12+6]) ^ ( R3[8+6] & R3[13+6]) ^ ( R3[13+6] & R3[15+6]) ^ ( R3[2+6] & R3[12+6] & R3[13+6]) ^ ( R3[7+6] & R3[8+6] & R3[12+6]) ^ ( R3[7+6] & R3[8+6] & R3[14+6]) ^ ( R3[8+6] & R3[12+6] & R3[13+6]) ^ ( R3[2+6] & R3[7+6] & R3[12+6] & R3[13+6]) ^ ( R3[2+6] & R3[7+6] & R3[13+6] & R3[14+6]) ^ ( R3[4+6] & R3[11+6] & R3[12+6] & R3[24+6]) ^ ( R3[7+6] & R3[8+6] & R3[12+6] & R3[13+6]) ^ ( R3[7+6] & R3[8+6] & R3[13+6] & R3[14+6]) ^ ( R3[4+6] & R3[7+6] & R3[11+6] & R3[12+6] & R3[24+6]) ^ ( R3[4+6] & R3[7+6] & R3[11+6] & R3[14+6] & R3[24+6]);
	assign F4p7_ = R4[0+6] ^ R4[2+6] ^ R4[7+6] ^ R4[9+6] ^ R4[10+6] ^ R4[15+6] ^ R4[23+6] ^ R4[25+6] ^ F1p4 ^ ( R4[8+6] & R4[15+6]) ^ ( R4[12+6] & R4[16+6]) ^ ( R4[13+6] & R4[15+6]) ^ ( R4[13+6] & R4[25+6]) ^ ( R4[1+6] & R4[8+6] & R4[14+6]) ^ ( R4[1+6] & R4[8+6] & R4[18+6]) ^ ( R4[8+6] & R4[12+6] & R4[16+6]) ^ ( R4[8+6] & R4[14+6] & R4[18+6]) ^ ( R4[8+6] & R4[15+6] & R4[16+6]) ^ ( R4[8+6] & R4[15+6] & R4[17+6]) ^ ( R4[15+6] & R4[17+6] & R4[24+6]) ^ ( R4[1+6] & R4[8+6] & R4[14+6] & R4[17+6]) ^ ( R4[1+6] & R4[8+6] & R4[17+6] & R4[18+6]) ^ ( R4[1+6] & R4[14+6] & R4[17+6] & R4[24+6]) ^ ( R4[1+6] & R4[17+6] & R4[18+6] & R4[24+6]) ^ ( R4[8+6] & R4[12+6] & R4[16+6] & R4[17+6]) ^ ( R4[8+6] & R4[14+6] & R4[17+6] & R4[18+6]) ^ ( R4[8+6] & R4[15+6] & R4[16+6] & R4[17+6]) ^ ( R4[12+6] & R4[16+6] & R4[17+6] & R4[24+6]) ^ ( R4[14+6] & R4[17+6] & R4[18+6] & R4[24+6]) ^ ( R4[15+6] & R4[16+6] & R4[17+6] & R4[24+6]);
	
	assign F1p7 = (state == State_Load_IV)? F1p7_ ^ iv[0+6] : F1p7_;
	assign F2p7 = (state == State_Load_IV)? F2p7_ ^ iv[0+6] : F2p7_;
	assign F3p7 = (state == State_Load_IV)? F3p7_ ^ iv[0+6] : F3p7_;
	assign F4p7 = (state == State_Load_IV)? F4p7_ ^ iv[0+6] : F4p7_;
	
	//-----Feedback function of P8---------
	assign F1p8_ = R1[0+7] ^ R1[2+7] ^ R1[5+7] ^ R1[6+7] ^ R1[15+7] ^ R1[17+7] ^ R1[18+7] ^ R1[20+7] ^ F4p2 ^ (R1[8+7] & R1[18+7]) ^ (R1[8+7] & R1[20+7]) ^ (R1[12+7] & R1[21+7]) ^ (R1[14+7] & R1[19+7]) ^ (R1[17+7] & R1[21+7]) ^ ( R1[20+7] & R1[22+7]) ^ ( R1[4+7] & R1[12+7] & R1[22+7]) ^ ( R1[4+7] & R1[19+7] & R1[22+7]) ^ ( R1[7+7] & R1[20+7] & R1[21+7]) ^ ( R1[8+7] & R1[18+7] & R1[22+7]) ^ ( R1[8+7] & R1[20+7] & R1[22+7]) ^ ( R1[12+7] & R1[19+7] & R1[22+7]) ^ ( R1[20+7] & R1[21+7] & R1[22+7]) ^ ( R1[4+7] & R1[7+7] & R1[12+7] & R1[21+7]) ^ ( R1[4+7] & R1[7+7] & R1[19+7] & R1[21+7]) ^ ( R1[4+7] & R1[12+7] & R1[21+7] & R1[22+7]) ^ ( R1[4+7] & R1[19+7] & R1[21+7] & R1[22+7]) ^ ( R1[7+7] & R1[8+7] & R1[18+7] & R1[21+7]) ^ ( R1[7+7] & R1[8+7] & R1[20+7] & R1[21+7]) ^ ( R1[7+7] & R1[12+7] & R1[19+7] & R1[21+7]) ^ ( R1[8+7] & R1[18+7] & R1[21+7] & R1[22+7]) ^ ( R1[8+7] & R1[20+7] & R1[21+7] & R1[22+7]) ^ ( R1[12+7] & R1[19+7] & R1[21+7] & R1[22+7]);
	assign F2p8_ = R2[0+7] ^ R2[3+7] ^ R2[17+7] ^ R2[22+7] ^ F3p4  ^ ( R2[2+7] & R2[13+7]) ^ ( R2[5+7] & R2[19+7]) ^ ( R2[7+7] & R2[19+7]) ^ ( R2[8+7] & R2[12+7]) ^ ( R2[8+7] & R2[13+7]) ^ ( R2[13+7] & R2[15+7]) ^ ( R2[2+7] & R2[12+7] & R2[13+7]) ^ ( R2[7+7] & R2[8+7] & R2[12+7]) ^ ( R2[7+7] & R2[8+7] & R2[14+7]) ^ ( R2[8+7] & R2[12+7] & R2[13+7]) ^ ( R2[2+7] & R2[7+7] & R2[12+7] & R2[13+7]) ^ ( R2[2+7] & R2[7+7] & R2[13+7] & R2[14+7]) ^ ( R2[4+7] & R2[11+7] & R2[12+7] & R2[24+7]) ^ ( R2[7+7] & R2[8+7] & R2[12+7] & R2[13+7]) ^ ( R2[7+7] & R2[8+7] & R2[13+7] & R2[14+7]) ^ ( R2[4+7] & R2[7+7] & R2[11+7] & R2[12+7] & R2[24+7]) ^ ( R2[4+7] & R2[7+7] & R2[11+7] & R2[14+7] & R2[24+7]);
	assign F3p8_ = R3[0+7] ^ R3[3+7] ^ R3[17+7] ^ R3[22+7] ^ F4p4  ^ ( R3[2+7] & R3[13+7]) ^ ( R3[5+7] & R3[19+7]) ^ ( R3[7+7] & R3[19+7]) ^ ( R3[8+7] & R3[12+7]) ^ ( R3[8+7] & R3[13+7]) ^ ( R3[13+7] & R3[15+7]) ^ ( R3[2+7] & R3[12+7] & R3[13+7]) ^ ( R3[7+7] & R3[8+7] & R3[12+7]) ^ ( R3[7+7] & R3[8+7] & R3[14+7]) ^ ( R3[8+7] & R3[12+7] & R3[13+7]) ^ ( R3[2+7] & R3[7+7] & R3[12+7] & R3[13+7]) ^ ( R3[2+7] & R3[7+7] & R3[13+7] & R3[14+7]) ^ ( R3[4+7] & R3[11+7] & R3[12+7] & R3[24+7]) ^ ( R3[7+7] & R3[8+7] & R3[12+7] & R3[13+7]) ^ ( R3[7+7] & R3[8+7] & R3[13+7] & R3[14+7]) ^ ( R3[4+7] & R3[7+7] & R3[11+7] & R3[12+7] & R3[24+7]) ^ ( R3[4+7] & R3[7+7] & R3[11+7] & R3[14+7] & R3[24+7]);
	assign F4p8_ = R4[0+7] ^ R4[2+7] ^ R4[7+7] ^ R4[9+7] ^ R4[10+7] ^ R4[15+7] ^ R4[23+7] ^ R4[25+7] ^ F4p5 ^ ( R4[8+7] & R4[15+7]) ^ ( R4[12+7] & R4[16+7]) ^ ( R4[13+7] & R4[15+7]) ^ ( R4[13+7] & R4[25+7]) ^ ( R4[1+7] & R4[8+7] & R4[14+7]) ^ ( R4[1+7] & R4[8+7] & R4[18+7]) ^ ( R4[8+7] & R4[12+7] & R4[16+7]) ^ ( R4[8+7] & R4[14+7] & R4[18+7]) ^ ( R4[8+7] & R4[15+7] & R4[16+7]) ^ ( R4[8+7] & R4[15+7] & R4[17+7]) ^ ( R4[15+7] & R4[17+7] & R4[24+7]) ^ ( R4[1+7] & R4[8+7] & R4[14+7] & R4[17+7]) ^ ( R4[1+7] & R4[8+7] & R4[17+7] & R4[18+7]) ^ ( R4[1+7] & R4[14+7] & R4[17+7] & R4[24+7]) ^ ( R4[1+7] & R4[17+7] & R4[18+7] & R4[24+7]) ^ ( R4[8+7] & R4[12+7] & R4[16+7] & R4[17+7]) ^ ( R4[8+7] & R4[14+7] & R4[17+7] & R4[18+7]) ^ ( R4[8+7] & R4[15+7] & R4[16+7] & R4[17+7]) ^ ( R4[12+7] & R4[16+7] & R4[17+7] & R4[24+7]) ^ ( R4[14+7] & R4[17+7] & R4[18+7] & R4[24+7]) ^ ( R4[15+7] & R4[16+7] & R4[17+7] & R4[24+7]);
	
	assign F1p8 = (state == State_Load_IV)? F1p8_ ^ iv[0+7] : F1p8_;
	assign F2p8 = (state == State_Load_IV)? F2p8_ ^ iv[0+7] : F2p8_;
	assign F3p8 = (state == State_Load_IV)? F3p8_ ^ iv[0+7] : F3p8_;
	assign F4p8 = (state == State_Load_IV)? F4p8_ ^ iv[0+7] : F4p8_;

endmodule 